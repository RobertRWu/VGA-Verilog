//////////////////////////////////////////////////////////////////////////////////
// Engineer: Robert Wu
// Create Date: 07/11/2019
// Project Name: VGA
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module VGA_char(
    input rst,
    input [2:0] h_index,
    input [3:0] v_index,
    input [4:0] a_index, 
    output reg point
    );

    reg [127:0] font_rom[16:0];
    wire [127:0] character;

    always @(posedge rst)
    begin
        if(rst) begin
            font_rom[0]  = {8'h00, 8'h00, 8'h3E, 8'h63, 8'h63, 8'h63, 8'h6B, 8'h6B, 8'h63, 8'h63, 8'h63, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00}; // 0
            font_rom[1]  = {8'h00, 8'h00, 8'h0C, 8'h1C, 8'h3C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00}; // 1
            font_rom[2]  = {8'h00, 8'h00, 8'h3E, 8'h63, 8'h03, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h61, 8'h63, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h00}; // 2
            font_rom[3]  = {8'h00, 8'h00, 8'h3E, 8'h63, 8'h03, 8'h03, 8'h1E, 8'h03, 8'h03, 8'h03, 8'h63, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00}; // 3
            font_rom[4]  = {8'h00, 8'h00, 8'h06, 8'h0E, 8'h1E, 8'h36, 8'h66, 8'h66, 8'h7F, 8'h06, 8'h06, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00}; // 4
            font_rom[5]  = {8'h00, 8'h00, 8'h7F, 8'h60, 8'h60, 8'h60, 8'h7E, 8'h03, 8'h03, 8'h63, 8'h73, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00}; // 5
            font_rom[6]  = {8'h00, 8'h00, 8'h1C, 8'h30, 8'h60, 8'h60, 8'h7E, 8'h63, 8'h63, 8'h63, 8'h63, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00}; // 6
            font_rom[7]  = {8'h00, 8'h00, 8'h7F, 8'h63, 8'h03, 8'h06, 8'h06, 8'h0C, 8'h0C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00}; // 7
            font_rom[8]  = {8'h00, 8'h00, 8'h3E, 8'h63, 8'h63, 8'h63, 8'h3E, 8'h63, 8'h63, 8'h63, 8'h63, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00}; // 8
            font_rom[9]  = {8'h00, 8'h00, 8'h3E, 8'h63, 8'h63, 8'h63, 8'h63, 8'h3F, 8'h03, 8'h03, 8'h06, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00}; // 9
            font_rom[10] = {8'h00, 8'h00, 8'h08, 8'h1C, 8'h36, 8'h63, 8'h63, 8'h63, 8'h7F, 8'h63, 8'h63, 8'h63, 8'h00, 8'h00, 8'h00, 8'h00}; // A
            font_rom[11] = {8'h00, 8'h00, 8'h7E, 8'h33, 8'h33, 8'h33, 8'h3E, 8'h33, 8'h33, 8'h33, 8'h33, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00}; // B
            font_rom[12] = {8'h00, 8'h00, 8'h1E, 8'h33, 8'h61, 8'h60, 8'h60, 8'h60, 8'h60, 8'h61, 8'h33, 8'h1E, 8'h00, 8'h00, 8'h00, 8'h00}; // C
            font_rom[13] = {8'h00, 8'h00, 8'h7C, 8'h36, 8'h33, 8'h33, 8'h33, 8'h33, 8'h33, 8'h33, 8'h36, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00}; // D
            font_rom[14] = {8'h00, 8'h00, 8'h7F, 8'h33, 8'h31, 8'h34, 8'h3C, 8'h34, 8'h30, 8'h31, 8'h33, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h00}; // E
            font_rom[15] = {8'h00, 8'h00, 8'h7F, 8'h33, 8'h31, 8'h34, 8'h3C, 8'h34, 8'h30, 8'h30, 8'h30, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00}; // F
            font_rom[16] = {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}; // space
        end
    end

    assign character = font_rom[a_index];   //alphabet index
    
    always @(*)
    begin
        point <= character[127 - (8*v_index + h_index)]; 
    end
    
endmodule
